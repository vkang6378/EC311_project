module word (
    input wire [4:0] rom_addr,
    output wire [0:127] M
);

    reg [0:127] rom[0:31];
    parameter data = {
    128'h00000000000000000000000000000000, 
    128'h00000000000000000000000000000000, 
    128'h003007000000e00001801e000003c000, 
    128'h1e3c0f800000f00001e01f000003e000, 
    128'h0f1e0f000000f70003e01e000003c018, 
    128'h0f9f0e000000f7c003c01e000003c03c, 
    128'h078f1e180018f3e007801e187ffffffe, 
    128'h078e1c3c003cf1f007801e3c3803c000, 
    128'h03c7dffe7ffef0f0070ffffe0003c000, 
    128'h00fff800383cf0780e3f1e000003c000, 
    128'h71fc38380038703c0e3c1e000703c1e0, 
    128'h7d9c7ffc00787ffe1c781e0007ffffe0, 
    128'h3d9c7e7c307fffc03cf01e000783c1c0, 
    128'h1f9cc0f03c7ff8607ff01e300783c1c0, 
    128'h1f9fe3e01e7078703fe01e780783c1c0, 
    128'h031de3c00ff078f83bc7fffc0783c1c0, 
    128'h073dc3c007f038f8038380000783c1c0, 
    128'h073dc3c003e039f00700000007ffffc0, 
    128'h0739c3dc01e03fe00e0f8070078fe1c0, 
    128'h0e39fffe01f03fc01ffffff8079ff1c0, 
    128'h7e39fbc003f83f803fe3c078071ff800, 
    128'h7e39c3c003f81f0c3f03c070003ffc00, 
    128'h3e71c3c007fc1e0c1c03c070007bde00, 
    128'h1e71c3c0073c3f0c0007c07000f3df00, 
    128'h1ef1c3c00e1c7f8c007fc07001f3cf80, 
    128'h1ee3c3c01e1df7cc07fbc07003c3c7e0, 
    128'h1de383c01c03e3fc7fc3c0700783c3fe, 
    128'h1dff83c0380783fc7f03fff01f03c1fe, 
    128'h1f9f9fc0701f01fc3c03c0703c03c078, 
    128'h070f0780e03c007e3003c0707803c030, 
    128'h060c03800030001e0003c07000038000, 
    128'h00000000000000000000000000000000
    };

    integer i;
    initial begin   //初始化，将data的数值输入到rom中
        for (i = 0;i < 32;i = i +1) 
            rom[i] = data[(4095-128*i)-:128];
    end

    assign M= rom[rom_addr];
endmodule